module Design1TB